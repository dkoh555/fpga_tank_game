library IEEE;
use IEEE.std_logic_1164.all;

--Additional standard or custom libraries go here
package tank_const is
	constant SCREEN_WIDTH : natural := 640;
	constant SCREEN_HEIGHT : natural := 480;
	constant TANK_WIDTH : natural := 80;
	constant TANK_HEIGHT : natural := 40;
	constant BULLET_SIZE : natural := 10;

end package tank_const;

package body tank_const is

end package body tank_const;