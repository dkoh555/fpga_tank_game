library IEEE;
use IEEE.std_logic_1164.all;

--Additional standard or custom libraries go here
package score_const is
	constant SCORE_WIDTH : natural := 2;
	constant WINNING_SCORE : natural := 3;
end package score_const;

package body score_const is

end package body score_const;